module transmitter_FSM(
    input logic baud_tick,
    output logic start, stop,
    output logic select
);


endmodule