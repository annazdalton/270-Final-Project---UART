`timescale 1ns / 1ps

module tb_transmitter_FSM();


endmodule