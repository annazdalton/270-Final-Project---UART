module transmitterMux(
    input logic piso_i, start, stop, parity_i,
    input logic [1:0] select,
    output logic tx_data_o
);


endmodule 